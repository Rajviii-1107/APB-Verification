`ifndef APB_DEFINES
`define APB_DEFINES

`define ADDR_WIDTH 32
`define DATA_WIDTH 32

`endif
